library verilog;
use verilog.vl_types.all;
entity question62 is
    port(
        L2              : out    vl_logic;
        Clock           : in     vl_logic;
        ResetLow        : in     vl_logic;
        L3              : out    vl_logic;
        L4              : out    vl_logic
    );
end question62;
