library verilog;
use verilog.vl_types.all;
entity question57_vlg_vec_tst is
end question57_vlg_vec_tst;
