library verilog;
use verilog.vl_types.all;
entity proj01 is
    port(
        C               : out    vl_logic;
        A               : in     vl_logic;
        B               : in     vl_logic
    );
end proj01;
