library verilog;
use verilog.vl_types.all;
entity question57_vlg_check_tst is
    port(
        out1            : in     vl_logic;
        out2            : in     vl_logic;
        out3            : in     vl_logic;
        out4            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end question57_vlg_check_tst;
