library verilog;
use verilog.vl_types.all;
entity Lab2 is
    port(
        D               : out    vl_logic;
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        SimpD           : out    vl_logic
    );
end Lab2;
