library verilog;
use verilog.vl_types.all;
entity question57 is
    port(
        out1            : out    vl_logic;
        clock           : in     vl_logic;
        out2            : out    vl_logic;
        out3            : out    vl_logic;
        out4            : out    vl_logic
    );
end question57;
