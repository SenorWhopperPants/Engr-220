library verilog;
use verilog.vl_types.all;
entity proj01_vlg_check_tst is
    port(
        C               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end proj01_vlg_check_tst;
