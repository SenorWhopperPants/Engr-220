library verilog;
use verilog.vl_types.all;
entity moore_state_machine_vlg_vec_tst is
end moore_state_machine_vlg_vec_tst;
