library verilog;
use verilog.vl_types.all;
entity proj01_vlg_vec_tst is
end proj01_vlg_vec_tst;
