library verilog;
use verilog.vl_types.all;
entity question62_vlg_vec_tst is
end question62_vlg_vec_tst;
