library verilog;
use verilog.vl_types.all;
entity question62_vlg_check_tst is
    port(
        L2              : in     vl_logic;
        L3              : in     vl_logic;
        L4              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end question62_vlg_check_tst;
